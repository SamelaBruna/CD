entity contadorModulo is
  port(A: in bit_vector(3 downto 0);
       bUD,Clr,load,en,Clock: in bit; 
       S: out bit_vector(3 downto 0)
       
       
    );
end contadorModulo;

architecture funcionamento of contadorModulo is

component JK is
     port (clk,J,K,P,C: IN BIT;
           q: OUT BIT
                   
     ); 
 end component; 

    signal inJK, logicPres,logicClr,outJK: bit_vector (3 downto 0);
    signal up,down: bit_vector(3 downto 0);   
    signal if10,if15: bit; 

 begin       

    logicPres(3)<=((not A(3)) or (not load) or Clr);
    logicPres(2)<=((not A(2)) or (not load) or Clr);
    logicPres(1)<=((not A(1)) or (not load) or Clr);
    logicPres(0)<=((not A(0)) or (not load) or Clr);


    logicClr(3)<=(not Clr) and ((load and A(3)) or (A(3) and not if10) or (not load and not if10));
    logicClr(2)<=(not Clr) and ((load and A(2)) or (A(2) and not if15) or (not load and not if15));
    logicClr(1)<=(not Clr) and ((load and A(1)) or (A(1) and not (if10 or if15)) or (not load and not (if10 or if15)));
    logicClr(0)<=(not Clr) and (not load or A(0));

    inJK(0)<=en;

    up(1)<=outJK(0) and not bUD;
    down(1)<=not outJK(0) and bUD;

    inJK(1)<=en and (up(1) or down(1));

    up(2)<=outJK(1) and up(1);
    down(2)<=not outJK(1) and down(1);

    inJK(2)<=en and (up(2) or down(2));

    up(3)<=outJK(2) and up(2);
    down(3)<=not outJK(2) and down(2);

    inJK(3)<=en and (up(3) or down(3));

   
    if10<=(outJK(3) and not outJK(2) and outJK(1) and not outJK(0)); --1010
    if15<=(outJK(3) and outJK(2) and outJK(1) and outJK(0)); --1111


    JK3: JK port map (
        clk => Clock,
        J=> inJK(3),
        K => inJK(3),
        P => logicPres(3),
        C=> logicClr(3),
        q => outJK(3)
        
    );

    JK2: JK port map (
        clk => Clock,
        J=> inJK(2),
        K => inJK(2),
        P => logicPres(2),
        C=> logicClr(2),
        q => outJK(2)
        
    );

    JK1: JK port map (
        clk => Clock,
        J=> inJK(1),
        K => inJK(1),
        P => logicPres(1),
        C=> logicClr(1),
        q => outJK(1)
        
    );

    JK0: JK port map (
        clk => Clock,
        J=> inJK(0),
        K => inJK(0),
        P => logicPres(0),
        C=> logicClr(0),
        q => outJK(0)
        
    );
          
    S <= outJK;

end funcionamento;
